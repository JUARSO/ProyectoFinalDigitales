module pruebaConexionRam(input [7:0] ram_Out [64:0]);



		



endmodule
