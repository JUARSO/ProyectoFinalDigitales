module pruebaConexionRam(input [7:0] ram_Out [64:0]);



always @(*)

		$display("%p",ram_Out[0]);


endmodule
