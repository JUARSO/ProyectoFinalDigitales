module modulo_PC(input logic clk, reset, output logic[31:0] pc);

	logic [31:0] pc_next;
	

	
	clk_pc #(32)  clkPc(clk, reset,pc_next,pc);
	sum_pc #(32) sumPC(pc,32'b100,pc_next);
	
	endmodule
	